`timescale 1ns/1ns

module ADD_1(
	input [31:0]A,
	output [31:0]result
);

assign result = A+4;

endmodule
